`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:   22:30:52 01/30/2011
// Design Name:   MiniAlu
// Module Name:   D:/Proyecto/RTL/Dev/MiniALU/TestBench.v
// Project Name:  MiniALU
// Target Device:
// Tool versions:
// Description:
//
// Verilog Test Fixture created by ISE for module: MiniAlu
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
////////////////////////////////////////////////////////////////////////////////

module TestBench(input clk);

// Inputs
reg Clock;
reg Reset;
wire rWrite;
wire [7: 0] rData;
wire wReady;


// Outputs
wire oLCD_Enabled;
wire oLCD_RegisterSelect;
wire oLCD_StrataFlashControl;
wire oLCD_ReadWrite;
wire [3: 0] oLCD_Data;
wire [7: 0] oLed;


// Instantiate the Unit Under Test (UUT)
MiniAlu uut (
          .Clock(Clock),
          .Reset(Reset),
          .oLed(oLed),
          .oLCD_Enabled(oLCD_Enabled),
          .oLCD_RegisterSelect(oLCD_RegisterSelect),
          .oLCD_StrataFlashControl(oLCD_StrataFlashContro),
          .oLCD_ReadWrite(oLCD_StrataFlashContro),
          .oLCD_Data(oLCD_Data)
        );

always
  begin
    #5 Clock = ! Clock;

  end

initial
  begin
    // Initialize Inputs
    Clock = 0;
    Reset = 0;

    // Wait 100 ns for global reset to finish
    #100;
    Reset = 1;
    #50
     Reset = 0;

    // Add stimulus here

  end

endmodule
