
`timescale 1ns / 1ps
`include "Defintions.v"
`include "Maquina_Estados.v"


module MiniAlu
       (
         input wire Clock,
         input wire Reset,
         output wire [7: 0] oLed,
         output wire wReady,
         output wire oLCD_Enabled,
         output wire oLCD_RegisterSelect,  //0=Command, 1=Data
         output wire oLCD_StrataFlashControl,
         output wire oLCD_ReadWrite,
         output wire [3: 0] oLCD_Data,
         input wire wWrite


       );

wire [15: 0] wIP, wIP_temp;
reg rWriteEnable, rBranchTaken;
wire [27: 0] wInstruction;
wire [3: 0] wOperation;
reg signed [15: 0] rResult, rResultHI; //Con signo
reg signed [31: 0] rResultTotal;
wire [7: 0] wSourceAddr0, wSourceAddr1, wDestination;
wire signed [15: 0] wSourceData0, wSourceData1, wIPInitialValue, wImmediateValue; //Con signo
wire [7: 0] rData;
wire rWrite;


ROM InstructionRom
    (
      .iAddress( wIP ),
      .oInstruction( wInstruction )
    );

RAM_DUAL_READ_PORT DataRam
                   (
                     .Clock( Clock ),
                     .iWriteEnable( rWriteEnable ),
                     .iReadAddress0( wInstruction[7: 0] ),
                     .iReadAddress1( wInstruction[15: 8] ),
                     .iWriteAddress( wDestination ),
                     .iDataIn( rResult ),
                     .oDataOut0( wSourceData0 ),
                     .oDataOut1( wSourceData1 )
                   );

assign wIPInitialValue = (Reset) ? 8'b0 : wDestination;
UPCOUNTER_POSEDGE IP
                  (
                    .Clock( Clock ),
                    .Reset( Reset | rBranchTaken ),
                    .Initial( wIPInitialValue + 16'd1 ),
                    .Enable( 1'b1 ),
                    .Q( wIP_temp )
                  );
assign wIP = (rBranchTaken) ? wIPInitialValue : wIP_temp;

FFD_POSEDGE_SYNCRONOUS_RESET # ( 4 ) FFD1
                             (
                               .Clock(Clock),
                               .Reset(Reset),
                               .Enable(1'b1),
                               .D(wInstruction[27: 24]),
                               .Q(wOperation)
                             );

FFD_POSEDGE_SYNCRONOUS_RESET # ( 8 ) FFD2
                             (
                               .Clock(Clock),
                               .Reset(Reset),
                               .Enable(1'b1),
                               .D(wInstruction[7: 0]),
                               .Q(wSourceAddr0)
                             );

FFD_POSEDGE_SYNCRONOUS_RESET # ( 8 ) FFD3
                             (
                               .Clock(Clock),
                               .Reset(Reset),
                               .Enable(1'b1),
                               .D(wInstruction[15: 8]),
                               .Q(wSourceAddr1)
                             );

FFD_POSEDGE_SYNCRONOUS_RESET # ( 8 ) FFD4
                             (
                               .Clock(Clock),
                               .Reset(Reset),
                               .Enable(1'b1),
                               .D(wInstruction[23: 16]),
                               .Q(wDestination)
                             );


reg rFFLedEN;
FFD_POSEDGE_SYNCRONOUS_RESET # ( 8 ) FF_LEDS
                             (
                               .Clock(Clock),
                               .Reset(Reset),
                               .Enable( rFFLedEN ),
                               .D( wSourceData1[7: 0] ),
                               .Q( oLed )
                             );

assign wImmediateValue = {wSourceAddr1, wSourceAddr0};

//Se instancia un ARRAY_MULT_GEN
// ARRAY_MULT_GEN # ( 16 ) arr_mul_gen
// (
//   .iMulA(wSourceData0),
//   .iMulB(wSourceData1),
//   .oMulR(wArrayMultGen)
// );

Module_LCD_Control LCD (
                     .Clock ( Clock ) ,
                     .Reset ( Reset ) ,
                     .wWrite ( rWrite ) ,
                     .wData ( rData ) ,
                     .wReady ( wReady ) ,
                     .oLCD_Enabled ( oLCD_Enabled ) ,
                     .oLCD_RegisterSelect ( oLCD_RegisterSelect ) ,  //0=Command, 1=Data
                     .oLCD_StrataFlashControl ( oLCD_StrataFlashControl ) ,
                     .oLCD_ReadWrite ( oLCD_ReadWrite ) ,
                     .oLCD_Data(oLCD_Data)
                   );



always @ ( * )
  begin
    case (wOperation)
      //-------------------------------------
      `NOP:
        begin
          rFFLedEN <= 1'b0;
          rBranchTaken <= 1'b0;
          rWriteEnable <= 1'b0;
          rResult <= 0;
        end

      //-------------------------------------
      `ADD:
        begin
          rFFLedEN <= 1'b0;
          rBranchTaken <= 1'b0;
          rWriteEnable <= 1'b1;
          rResult <= wSourceData1 + wSourceData0;
        end

      //-------------------------------------
      `SUB:
        begin
          rFFLedEN <= 1'b0;
          rBranchTaken <= 1'b0;
          rWriteEnable <= 1'b1;
          rResult <= wSourceData1 - wSourceData0;
        end

      //-------------------------------------
      `STO:
        begin
          rFFLedEN <= 1'b0;
          rWriteEnable <= 1'b1;
          rBranchTaken <= 1'b0;
          rResult <= wImmediateValue;
        end

      //-------------------------------------
      `BLE:
        begin
          rFFLedEN <= 1'b0;
          rWriteEnable <= 1'b0;
          rResult <= 0;

          if (wSourceData1 <= wSourceData0 )
            rBranchTaken <= 1'b1;
          else
            rBranchTaken <= 1'b0;

        end

      //-------------------------------------
      `JMP:
        begin
          rFFLedEN <= 1'b0;
          rWriteEnable <= 1'b0;
          rResult <= 0;
          rBranchTaken <= 1'b1;
        end

      //-------------------------------------
      `LED:
        begin
          rFFLedEN <= 1'b1;
          rWriteEnable <= 1'b0;
          rResult <= 0;
          rBranchTaken <= 1'b0;
        end

      //-------------------------------------
      //-------------------------------------
      `SMUL:
        begin
          rFFLedEN <= 1'b0;
          rBranchTaken <= 1'b0;
          rWriteEnable <= 1'b1;
          {rResultHI, rResult} <= wSourceData1 * wSourceData0;
          rResultTotal <= {rResultHI, rResult};
          //		rResult <= wSourceData1 * wSourceData0;
        end

      //-------------------------------------
      // `IMUL:
      // begin
      // 	rFFLedEN     <= 1'b0;
      // 	rBranchTaken <= 1'b0;
      // 	rWriteEnable <= 1'b1;
      // 	{rResultHI,rResult} <= wArrayMultGen;
      // 	rResultTotal <= {rResultHI,rResult};
      // end
      //-------------------------------------
      default:
        begin
          rFFLedEN <= 1'b1;
          rWriteEnable <= 1'b0;
          rResult <= 0;
          rBranchTaken <= 1'b0;
        end

      //-------------------------------------
    endcase
  end


endmodule
